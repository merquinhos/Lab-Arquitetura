// Módulo da Memória de Instruções usando um decodificador com 'case'
module instruction_memory_case (
    input  logic [31:0] a,   // Entrada de Endereço (do PC)
    output logic [31:0] rd  // Saída de Instrução (para o datapath)
);

    always_comb begin
        // obter o endereço da palavra (dividindo por 4).
        case (a[31:2])
				32'h00: rd = 32'h00700093; 
				32'h01: rd = 32'h00300193; 
				32'h02: rd = 32'hfff00113;  
				32'h03: rd = 32'h00110113;  
				32'h04: rd = 32'h003123b3; 
				32'h05: rd = 32'hfe208ae3; 
				32'h06: rd = 32'hfe000ae3; 
            
            default: rd = 32'h00000000;
        endcase
    end

endmodule


