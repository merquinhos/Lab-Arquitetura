// Code your design here
//porta xor 2x1
module xor2x1 (input logic a, b, output logic out);
  assign out = a^b;
  
endmodule

